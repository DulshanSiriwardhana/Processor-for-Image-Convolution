`timescale 1ns / 1ps
module control_unit(
	input clk,
	input enable,
	input Z_flag,
	input [5:0] addr,
	input [5:0] MBRU,
	output reg [37:0] control_signal,
	output finish
);

reg start = 1'b0;

reg [37:0] ROM[0:60];

reg check = 1'b0;

assign finish = check ;

// parameters
parameter FETCH2 = 6'd1;

parameter JUMPNZ = 6'd47;
parameter JUMPZ = 6'd52;

parameter JMPNZ1 = 6'd48;
parameter JMPNZY1 = 6'd49;

parameter JMPZN1 = 6'd53;
parameter JMPZY1 = 6'd54;
parameter JMPZY2 = 6'd55;

parameter NOP = 6'd46;


initial
	begin
		control_signal =38'b000000_0000_0000000000000000000_000_0_00000;
	end


always@ ( posedge enable )
	start = 1'b1;

always@(posedge clk)
	begin
		case(control_signal[37:32])
		FETCH2:
			begin
			control_signal = {MBRU, ROM[FETCH2][31:0]};
			end
		JUMPNZ:
			begin
				if (Z_flag == 1'b0)
					control_signal = {JMPNZ1, ROM[JMPNZ1][31:0]};
				else if (Z_flag == 1'b1)
					control_signal = {JMPZY1, ROM[JMPZY1][31:0]};
			end
		JUMPZ:
			begin
				if (Z_flag == 1'b0)
					control_signal = {JMPZN1, ROM[JMPZN1][31:0]};
				else if (Z_flag == 1'b1)
				 	control_signal = {JMPZY1, ROM[JMPZY1][31:0]};
			end
		
		NOP: 
			check = 1'b1;
	default : control_signal = ROM[addr];
	endcase
end

initial
begin

ROM[0] = 38'b000001_0000_0000000000000000000_100_0_00000; //FETCH1
ROM[1] = 38'bxxxxxx_0000_0000000000000000000_000_1_00000; //FETCH2
ROM[2] = 38'b000000_1001_0000000000000000001_000_0_00000; //CLAC
ROM[3] = 38'b000000_0101_1000000000000000000_000_0_00000; //MVACMAR
ROM[4] = 38'b000101_0000_0000000000000000000_010_0_00000; //LDAC1
//ROM[5] = 38'b000000_0110_0000000000000000001_000_0_00001; //LDAC2

//
ROM[5] = 38'b000000_0110_0000000000000000001_000_0_00001; //LDAC2
ROM[5] = 38'b000000_0110_0000000000000000001_000_0_00001; //LDAC2

ROM[6] = 38'b000000_0101_0001000000000000000_000_0_00000; //MVACK0
ROM[7] = 38'b000000_0111_0000000000000000001_000_0_00000; //INAC
ROM[8] = 38'b000000_0101_0000000000000000010_000_0_00000; //MVACI
ROM[9] = 38'b000000_0101_0000100000000000000_000_0_00000; //MVACK1
ROM[10] = 38'b000000_0110_0000000000000000001_000_0_10000; //MVIAC
ROM[11] = 38'b000000_0101_0000010000000000000_000_0_00000; //MVACK2
ROM[12] = 38'b000000_0101_0000001000000000000_000_0_00000; //MVACK3
ROM[13] = 38'b000000_0101_0000000100000000000_000_0_00000; //MVACK4
ROM[14] = 38'b000000_0101_0000000010000000000_000_0_00000; //MVACK5
ROM[15] = 38'b000000_0101_0000000001000000000_000_0_00000; //MVACK6
ROM[16] = 38'b000000_0101_0000000000100000000_000_0_00000; //MVACK7
ROM[17] = 38'b000000_0101_0000000000010000000_000_0_00000; //MVACK8
ROM[18] = 38'b000000_0101_0000000000001000000_000_0_00000; //MVACP1
ROM[19] = 38'b000000_0110_0000000000000000010_000_0_10001; //LDII
//
//ROM[19] = 38'b000000_0001_0000000000000001000_000_0_10001; //LDII
//

//ROM[57] = 38'b000000_0101_0000000000000000010_000_0_00000; //LDII    MVACI
ROM[20] = 38'b000000_0101_0000000000000100000_000_0_00000; //MVACP2
//ROM[21] = 38'b000000_0001_0000000000000000001_000_0_10000; //ADDI
//
ROM[21] = 38'b111100_0001_0000000000000000000_000_0_10000; //ADDI
ROM[60] = 38'b000000_0000_0000000000000000001_000_0_00000; //ADDI

ROM[22] = 38'b000000_0101_0000000000000010000_000_0_00000; //MVACP3
ROM[23] = 38'b000000_0110_0000000000000001000_000_0_10001; //LDIDP
ROM[24] = 38'b000000_0101_0000000000000000100_000_0_00000; //MVACCV
ROM[25] = 38'b000000_0110_0000000000000000001_000_0_01011; //MVP1AC
ROM[26] = 38'b000000_0011_0000000000000000001_000_0_00010; //MULK0
ROM[27] = 38'b000000_0110_0000000000000000001_000_0_01100; //MVP2AC
ROM[28] = 38'b000000_0011_0000000000000000001_000_0_00101; //MULK3
ROM[29] = 38'b000000_0001_0000000000000000001_000_0_01111; //ADDCV
ROM[30] = 38'b000000_0011_0000000000000000001_000_0_01000; //MULK6
ROM[31] = 38'b000000_0011_0000000000000000001_000_0_00011; //MULK1
ROM[32] = 38'b000000_0011_0000000000000000001_000_0_00110; //MULK4
ROM[33] = 38'b000000_0110_0000000000000000001_000_0_01101; //MVP3AC
ROM[34] = 38'b000000_0011_0000000000000000001_000_0_01001; //MULK7
ROM[35] = 38'b000000_0011_0000000000000000001_000_0_00100; //MULK2
ROM[36] = 38'b000000_0011_0000000000000000001_000_0_00111; //MULK5
ROM[37] = 38'b000000_0011_0000000000000000001_000_0_01010; //MULK8
ROM[38] = 38'b000000_0110_0000000000000000001_000_0_01110; //MVDPAC
ROM[39] = 38'b000000_0101_0000000000000000100_000_0_00000; //MVCVAC
ROM[40] = 38'b000000_0100_0000000000000000001_000_0_00000; //MOD30
ROM[41] = 38'b101010_0101_0100000000000000000_000_0_00000; //STAC1
ROM[42] = 38'b000000_0000_0000000000000000000_001_0_00001; //STAC2 // check again
ROM[43] = 38'b000000_0110_0000000000000000010_000_0_10001; //MVII
//ROM[44] = 38'b000000_0010_0000000000000000001_000_0_10000; //SUBI
//ROM[44] = 38'b111010_0000_0000000000000000000_000_0_10000; //SUBI
//
ROM[44] = 38'b111010_0000_0000000000000000000_000_0_10000; //SUBI
ROM[58] = 38'b000000_0010_0000000000000000001_000_0_00000; //SUBI

ROM[45] = 38'b000000_0101_0000000000000001000_000_0_00000; //MVACDP
ROM[46] = 38'b000000_0000_0000000000000000000_000_0_00000; //NOP
ROM[47] = 38'bxxxxxx_0000_0000000000000000000_000_0_00000; //JUMPNZ
ROM[48] = 38'b000000_0000_0000000000000000000_000_0_00000; //JMPNZN1 Z = 0
//ROM[49] = 38'b110010_0110_0000000000000000001_100_0_10001; //JMPNZY1 Z = 1
//ROM[49] = 38'b111001_0000_0000000000000000000_000_0_10001; //JMPNZY1 Z = 1
ROM[49] = 38'b000000_0110_0000000000000000001_000_0_10001; //JMPNZY1 Z = 1


ROM[50] = 38'b110011_0101_0010000000000000001_000_0_00000; //JMPNZY2
ROM[51] = 38'b000000_0000_0000000000000000001_000_0_00000; //JMPNZY3
ROM[52] = 38'bxxxxxx_0000_0000000000000000000_000_0_00000; //JUMPZ
ROM[53] = 38'b000000_0000_0000000000000000000_000_0_00000; //JMPZN1 Z = 0
//ROM[54] = 38'b110111_0110_0000000000000000001_100_0_10001; //JMPZY1 Z = 1
 
// - ROM[54] = 38'b000000_0110_0000000000000000001_000_0_10001; //JMPZY1 Z = 1
ROM[54] = 38'b110111_0110_0000000000000000001_000_0_10001; //JMPZY1 Z = 1

ROM[55] = 38'b111000_0101_0010000000000000000_000_0_00000; //JMPZY2
ROM[56] = 38'b111001_0000_0000000000000000000_000_0_00000; //JMPZY2
ROM[57] = 38'b000000_1001_0000000000000000001_000_0_00000; //JMPZY2
ROM[59] = 38'b000000_1000_0000000000000000001_000_0_00000; //DECAC
//ROM[57] = 38'b111010_0110_0000000000000000000_000_0_00000; //LDII2
//ROM[58] = 38'b110010_0000_0000000000000000001_100_0_00000; //LDII2
//
//ROM[59] = 38'b110111_0110_0000000000000000001_100_0_00000; //LDII2
end

endmodule